magic
tech scmos
timestamp 1613729353
<< metal1 >>
rect -4 38 0 182
rect 512 42 519 182
rect 480 38 519 42
use oinverter  oinverter_1
array 0 15 -32 0 0 -110
timestamp 1613729060
transform -1 0 20 0 -1 172
box -12 -48 20 62
use oinverter  oinverter_0
array 0 14 32 0 0 110
timestamp 1613729060
transform 1 0 12 0 1 48
box -12 -48 20 62
<< end >>
