magic
tech scmos
timestamp 1613716236
<< nwell >>
rect -8 -5 17 62
<< ntransistor >>
rect 4 -33 6 -13
<< ptransistor >>
rect 4 1 6 51
<< ndiffusion >>
rect 3 -33 4 -13
rect 6 -33 7 -13
<< pdiffusion >>
rect 3 1 4 51
rect 6 1 7 51
<< ndcontact >>
rect -1 -33 3 -13
rect 7 -33 11 -13
<< pdcontact >>
rect -1 1 3 51
rect 7 1 11 51
<< polysilicon >>
rect 4 51 6 54
rect 4 -13 6 1
rect 4 -36 6 -33
<< polycontact >>
rect 0 -10 4 -6
<< metal1 >>
rect -8 58 17 62
rect -1 51 3 58
rect 7 -6 11 1
rect -10 -10 0 -6
rect 7 -10 20 -6
rect 7 -13 11 -10
rect -1 -44 3 -33
rect -8 -48 17 -44
<< labels >>
rlabel metal1 -8 -8 -8 -8 3 in
rlabel metal1 19 -8 19 -8 7 out
rlabel metal1 16 61 16 61 6 vdd
rlabel metal1 16 -46 16 -46 8 gnd
<< end >>
